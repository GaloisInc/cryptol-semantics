(* Copyright 2012-2015 by Adam Petcher.				*
 * Use of this source code is governed by the license described	*
 * in the LICENSE file at the root of the source tree.		*)
(* A top-level module that exports all of the common components of the framework. *)

Require Export otp.DistRules.
Require Export otp.Comp.
Require Export Arith.
Require Export otp.Fold.
Require Export otp.Rat.
Require Export otp.DistSem.
Require Export otp.StdNat.
Require Export otp.DistTacs.


Open Scope comp_scope.
Open Scope rat_scope.